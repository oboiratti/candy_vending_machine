library verilog;
use verilog.vl_types.all;
entity seven_seg_mux_tb is
end seven_seg_mux_tb;
