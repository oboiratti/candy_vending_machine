library verilog;
use verilog.vl_types.all;
entity key_map_tb is
end key_map_tb;
