library verilog;
use verilog.vl_types.all;
entity bcd_to_seven_seg_dec_tb is
end bcd_to_seven_seg_dec_tb;
